module MOD2 (A, B);

    input A;
    input B;

    wire A;
    wire B;
endmodule

// Some comment