

module top
(
    in1,
    in2,
    out1,
    out2,
);

    input in1;
    input [1:0]in2;
    output out1;
    output [1:0]out2;

endmodule

